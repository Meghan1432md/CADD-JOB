module c_tb;
    logic a, b, c, d;
    logic y, z;
    c uut (.a(a),.b(b),.c(c),.d(d),.y(y),.z(z));
    initial 
    begin
        a = 0; b = 0; c = 0; d = 0;
        #10 a = 1; b = 0; c = 0; d = 1;
        #10 a = 1; b = 1; c = 1; d = 1;
        #10 a = 0; b = 1; c = 0; d = 1;
        #10 a = 1; b = 1; c = 0; d = 0;
        #10 $finish;
    end
endmodule
